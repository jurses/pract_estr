module alu(output wire [3:0] R, output wire zero, carry, sign, input wire [3:0] A, B, input wire[1:0] AlUop, input wire L);
cal cal0(R[0], , A[0], B[1], );
endmodule
